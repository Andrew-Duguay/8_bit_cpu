library ieee;
use ieee.std_logic_1164.all;

entity ALU is
    port (
        z_flag   : out STD_LOGIC;
        n_flag   : out STD_LOGIC;
        v_flag   : out STD_LOGIC;
        c_flag   : out STD_LOGIC
    );
end entity ALU;

architecture rtl of ALU is
begin
    
end architecture rtl;    