library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

entity status_register_tb is
end entity status_register_tb;

architecture behavioral of status_register_tb is

begin

end architecture behavioral;
